//`define TEST_FILE "../sw/dmac_gpio_test.hex"
`define TEST_FILE "../FW/uart_test.hex"
`define VCD

